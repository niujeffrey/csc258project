module BrickBreaker();

endmodule

